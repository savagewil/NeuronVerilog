// neuron model
module backPropper(input wire [31:0] [31:0] bp_ds, input wire [32:0] [31:0] bp_w,
    input wire [63:0] bp_bp, input wire [31:0]  bp_tm, input wire [31:0]  bp_td,
    output wire [31:0] [31:0]  bp_bc, output reg [32:0] [31:0]  bp_wn);

    wire [31:0] test;
    backPropper_1 bp0(bp_ds[0], bp_w[0], bp_bp,  bp_tm,  bp_td,
         bp_bc[0],  bp_wn[0]);

    backPropper_1 bp1(bp_ds[1], bp_w[1], bp_bp,  bp_tm,  bp_td,
         bp_bc[1],  bp_wn[1]);

    backPropper_1 bp2(bp_ds[2], bp_w[2], bp_bp,  bp_tm,  bp_td,
         bp_bc[2],  bp_wn[2]);

    backPropper_1 bp3(bp_ds[3], bp_w[3], bp_bp,  bp_tm,  bp_td,
         bp_bc[3],  bp_wn[3]);

    backPropper_1 bp4(bp_ds[4], bp_w[4], bp_bp,  bp_tm,  bp_td,
         bp_bc[4],  bp_wn[4]);

    backPropper_1 bp5(bp_ds[5], bp_w[5], bp_bp,  bp_tm,  bp_td,
         bp_bc[5],  bp_wn[5]);

    backPropper_1 bp6(bp_ds[6], bp_w[6], bp_bp,  bp_tm,  bp_td,
         bp_bc[6],  bp_wn[6]);

    backPropper_1 bp7(bp_ds[7], bp_w[7], bp_bp,  bp_tm,  bp_td,
         bp_bc[7],  bp_wn[7]);

    backPropper_1 bp8(bp_ds[8], bp_w[8], bp_bp,  bp_tm,  bp_td,
         bp_bc[8],  bp_wn[8]);

    backPropper_1 bp9(bp_ds[9], bp_w[9], bp_bp,  bp_tm,  bp_td,
         bp_bc[9],  bp_wn[9]);

    backPropper_1 bp10(bp_ds[10], bp_w[10], bp_bp,  bp_tm,  bp_td,
         bp_bc[10],  bp_wn[10]);

    backPropper_1 bp11(bp_ds[11], bp_w[11], bp_bp,  bp_tm,  bp_td,
         bp_bc[11],  bp_wn[11]);

    backPropper_1 bp12(bp_ds[12], bp_w[12], bp_bp,  bp_tm,  bp_td,
         bp_bc[12],  bp_wn[12]);

    backPropper_1 bp13(bp_ds[13], bp_w[13], bp_bp,  bp_tm,  bp_td,
         bp_bc[13],  bp_wn[13]);

    backPropper_1 bp14(bp_ds[14], bp_w[14], bp_bp,  bp_tm,  bp_td,
         bp_bc[14],  bp_wn[14]);

    backPropper_1 bp15(bp_ds[15], bp_w[15], bp_bp,  bp_tm,  bp_td,
         bp_bc[15],  bp_wn[15]);

    backPropper_1 bp16(bp_ds[16], bp_w[16], bp_bp,  bp_tm,  bp_td,
         bp_bc[16],  bp_wn[16]);

    backPropper_1 bp17(bp_ds[17], bp_w[17], bp_bp,  bp_tm,  bp_td,
         bp_bc[17],  bp_wn[17]);

    backPropper_1 bp18(bp_ds[18], bp_w[18], bp_bp,  bp_tm,  bp_td,
         bp_bc[18],  bp_wn[18]);

    backPropper_1 bp19(bp_ds[19], bp_w[19], bp_bp,  bp_tm,  bp_td,
         bp_bc[19],  bp_wn[19]);

    backPropper_1 bp20(bp_ds[20], bp_w[20], bp_bp,  bp_tm,  bp_td,
         bp_bc[20],  bp_wn[20]);

    backPropper_1 bp21(bp_ds[21], bp_w[21], bp_bp,  bp_tm,  bp_td,
         bp_bc[21],  bp_wn[21]);

    backPropper_1 bp22(bp_ds[22], bp_w[22], bp_bp,  bp_tm,  bp_td,
         bp_bc[22],  bp_wn[22]);

    backPropper_1 bp23(bp_ds[23], bp_w[23], bp_bp,  bp_tm,  bp_td,
         bp_bc[23],  bp_wn[23]);

    backPropper_1 bp24(bp_ds[24], bp_w[24], bp_bp,  bp_tm,  bp_td,
         bp_bc[24],  bp_wn[24]);

    backPropper_1 bp25(bp_ds[25], bp_w[25], bp_bp,  bp_tm,  bp_td,
         bp_bc[25],  bp_wn[25]);

    backPropper_1 bp26(bp_ds[26], bp_w[26], bp_bp,  bp_tm,  bp_td,
         bp_bc[26],  bp_wn[26]);

    backPropper_1 bp27(bp_ds[27], bp_w[27], bp_bp,  bp_tm,  bp_td,
         bp_bc[27],  bp_wn[27]);

    backPropper_1 bp28(bp_ds[28], bp_w[28], bp_bp,  bp_tm,  bp_td,
         bp_bc[28],  bp_wn[28]);

    backPropper_1 bp29(bp_ds[29], bp_w[29], bp_bp,  bp_tm,  bp_td,
         bp_bc[29],  bp_wn[29]);

    backPropper_1 bp30(bp_ds[30], bp_w[30], bp_bp,  bp_tm,  bp_td,
         bp_bc[30],  bp_wn[30]);

    backPropper_1 bp31(bp_ds[31], bp_w[31], bp_bp,  bp_tm,  bp_td,
         bp_bc[31],  bp_wn[31]);

    backPropper_t bpthresh(bp_w[32], bp_bp,  bp_tm,  bp_td,
         bp_wn[32]);

endmodule: backPropper

