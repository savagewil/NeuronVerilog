module neuron(den1[31:0], den2[31:0], den3[31:0], den4[31:0], den5[31:0], den6[31:0], den7[31:0],
    den8[31:0], den9[31:0], den10[31:0], den11[31:0], den12[31:0], den13[31:0], den14[31:0],
    den15[31:0], den16[31:0], den17[31:0], den18[31:0], den19[31:0], den20[31:0], den21[31:0],
    den21[31:0], den23[31:0], den24[31:0], den25[31:0], den26[31:0], den27[31:0], den28[31:0],
    den29[31:0], den30[31:0], den31[31:0], den32[31:0], axon[31:0]);

    input den1, den2, den3, den4, den5, den6, den7, den8, den9, den10, den11, den12, den13, den14,
          den15, den16, den17, den18, den19, den20, den21, den21, den23, den24, den25, den26, den27,
          den28, den29, den30, den31, den32;
    output axon;


endmodule: neuron