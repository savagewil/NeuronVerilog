// neuron model
module backPropper(input wire [31:0] [31:0] dendrites, input wire [32:0] [31:0] weights,
    input wire [31:0] backprop, input wire [31:0] trainingMul, input wire [31:0] trainingDiv,
    output wire [31:0] [31:0] backpropChange, output wire [32:0] [31:0] weightNew);

    backPropper_1 bp0(dendrites[0], weights[0], backprop, trainingMul, trainingDiv,
        backpropChange[0], weightNew[0]);

    backPropper_1 bp1(dendrites[1], weights[1], backprop, trainingMul, trainingDiv,
        backpropChange[1], weightNew[1]);

    backPropper_1 bp2(dendrites[2], weights[2], backprop, trainingMul, trainingDiv,
        backpropChange[2], weightNew[2]);

    backPropper_1 bp3(dendrites[3], weights[3], backprop, trainingMul, trainingDiv,
        backpropChange[3], weightNew[3]);

    backPropper_1 bp4(dendrites[4], weights[4], backprop, trainingMul, trainingDiv,
        backpropChange[4], weightNew[4]);

    backPropper_1 bp5(dendrites[5], weights[5], backprop, trainingMul, trainingDiv,
        backpropChange[5], weightNew[5]);

    backPropper_1 bp6(dendrites[6], weights[6], backprop, trainingMul, trainingDiv,
        backpropChange[6], weightNew[6]);

    backPropper_1 bp7(dendrites[7], weights[7], backprop, trainingMul, trainingDiv,
        backpropChange[7], weightNew[7]);

    backPropper_1 bp8(dendrites[8], weights[8], backprop, trainingMul, trainingDiv,
        backpropChange[8], weightNew[8]);

    backPropper_1 bp9(dendrites[9], weights[9], backprop, trainingMul, trainingDiv,
        backpropChange[9], weightNew[9]);

    backPropper_1 bp10(dendrites[10], weights[10], backprop, trainingMul, trainingDiv,
        backpropChange[10], weightNew[10]);

    backPropper_1 bp11(dendrites[11], weights[11], backprop, trainingMul, trainingDiv,
        backpropChange[11], weightNew[11]);

    backPropper_1 bp12(dendrites[12], weights[12], backprop, trainingMul, trainingDiv,
        backpropChange[12], weightNew[12]);

    backPropper_1 bp13(dendrites[13], weights[13], backprop, trainingMul, trainingDiv,
        backpropChange[13], weightNew[13]);

    backPropper_1 bp14(dendrites[14], weights[14], backprop, trainingMul, trainingDiv,
        backpropChange[14], weightNew[14]);

    backPropper_1 bp15(dendrites[15], weights[15], backprop, trainingMul, trainingDiv,
        backpropChange[15], weightNew[15]);

    backPropper_1 bp16(dendrites[16], weights[16], backprop, trainingMul, trainingDiv,
        backpropChange[16], weightNew[16]);

    backPropper_1 bp17(dendrites[17], weights[17], backprop, trainingMul, trainingDiv,
        backpropChange[17], weightNew[17]);

    backPropper_1 bp18(dendrites[18], weights[18], backprop, trainingMul, trainingDiv,
        backpropChange[18], weightNew[18]);

    backPropper_1 bp19(dendrites[19], weights[19], backprop, trainingMul, trainingDiv,
        backpropChange[19], weightNew[19]);

    backPropper_1 bp20(dendrites[20], weights[20], backprop, trainingMul, trainingDiv,
        backpropChange[20], weightNew[20]);

    backPropper_1 bp21(dendrites[21], weights[21], backprop, trainingMul, trainingDiv,
        backpropChange[21], weightNew[21]);

    backPropper_1 bp22(dendrites[22], weights[22], backprop, trainingMul, trainingDiv,
        backpropChange[22], weightNew[22]);

    backPropper_1 bp23(dendrites[23], weights[23], backprop, trainingMul, trainingDiv,
        backpropChange[23], weightNew[23]);

    backPropper_1 bp24(dendrites[24], weights[24], backprop, trainingMul, trainingDiv,
        backpropChange[24], weightNew[24]);

    backPropper_1 bp25(dendrites[25], weights[25], backprop, trainingMul, trainingDiv,
        backpropChange[25], weightNew[25]);

    backPropper_1 bp26(dendrites[26], weights[26], backprop, trainingMul, trainingDiv,
        backpropChange[26], weightNew[26]);

    backPropper_1 bp27(dendrites[27], weights[27], backprop, trainingMul, trainingDiv,
        backpropChange[27], weightNew[27]);

    backPropper_1 bp28(dendrites[28], weights[28], backprop, trainingMul, trainingDiv,
        backpropChange[28], weightNew[28]);

    backPropper_1 bp29(dendrites[29], weights[29], backprop, trainingMul, trainingDiv,
        backpropChange[29], weightNew[29]);

    backPropper_1 bp30(dendrites[30], weights[30], backprop, trainingMul, trainingDiv,
        backpropChange[30], weightNew[30]);

    backPropper_1 bp31(dendrites[31], weights[31], backprop, trainingMul, trainingDiv,
        backpropChange[31], weightNew[31]);

    backPropper_t bpthresh(weights[32], backprop, trainingMul, trainingDiv,
        weightNew[32]);

endmodule: backPropper

