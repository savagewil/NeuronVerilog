module summer(
    input wire [32:0] [31:0] in,
    output reg [63:0]);
endmodule : summer