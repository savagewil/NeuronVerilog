// neuron model
module backPropper(input real bp_dendrites [31:0], input real bp_weights [32:0],
    input real bp_axon,
    input real bp_backprop,
    input real bp_training_ratio,
    output real bp_backprop_change [31:0],
    output real bp_weights_new [32:0]);

    backPropper_1 bp0(bp_dendrites[0],
        bp_weights[0],
        bp_axon,
        bp_backprop,
        bp_training_ratio,
        bp_backprop_change[0],
        bp_weights_new[0]);

    backPropper_1 bp1(bp_dendrites[1],
        bp_weights[1],
        bp_axon,
        bp_backprop,
        bp_training_ratio,
        bp_backprop_change[1],
        bp_weights_new[1]);

    backPropper_1 bp2(bp_dendrites[2],
        bp_weights[2],
        bp_axon,
        bp_backprop,
        bp_training_ratio,
        bp_backprop_change[2],
        bp_weights_new[2]);

    backPropper_1 bp3(bp_dendrites[3],
        bp_weights[3],
        bp_axon,
        bp_backprop,
        bp_training_ratio,
        bp_backprop_change[3],
        bp_weights_new[3]);

    backPropper_1 bp4(bp_dendrites[4],
        bp_weights[4],
        bp_axon,
        bp_backprop,
        bp_training_ratio,
        bp_backprop_change[4],
        bp_weights_new[4]);

    backPropper_1 bp5(bp_dendrites[5],
        bp_weights[5],
        bp_axon,
        bp_backprop,
        bp_training_ratio,
        bp_backprop_change[5],
        bp_weights_new[5]);

    backPropper_1 bp6(bp_dendrites[6],
        bp_weights[6],
        bp_axon,
        bp_backprop,
        bp_training_ratio,
        bp_backprop_change[6],
        bp_weights_new[6]);

    backPropper_1 bp7(bp_dendrites[7],
        bp_weights[7],
        bp_axon,
        bp_backprop,
        bp_training_ratio,
        bp_backprop_change[7],
        bp_weights_new[7]);

    backPropper_1 bp8(bp_dendrites[8],
        bp_weights[8],
        bp_axon,
        bp_backprop,
        bp_training_ratio,
        bp_backprop_change[8],
        bp_weights_new[8]);

    backPropper_1 bp9(bp_dendrites[9],
        bp_weights[9],
        bp_axon,
        bp_backprop,
        bp_training_ratio,
        bp_backprop_change[9],
        bp_weights_new[9]);

    backPropper_1 bp10(bp_dendrites[10],
        bp_weights[10],
        bp_axon,
        bp_backprop,
        bp_training_ratio,
        bp_backprop_change[10],
        bp_weights_new[10]);

    backPropper_1 bp11(bp_dendrites[11],
        bp_weights[11],
        bp_axon,
        bp_backprop,
        bp_training_ratio,
        bp_backprop_change[11],
        bp_weights_new[11]);

    backPropper_1 bp12(bp_dendrites[12],
        bp_weights[12],
        bp_axon,
        bp_backprop,
        bp_training_ratio,
        bp_backprop_change[12],
        bp_weights_new[12]);

    backPropper_1 bp13(bp_dendrites[13],
        bp_weights[13],
        bp_axon,
        bp_backprop,
        bp_training_ratio,
        bp_backprop_change[13],
        bp_weights_new[13]);

    backPropper_1 bp14(bp_dendrites[14],
        bp_weights[14],
        bp_axon,
        bp_backprop,
        bp_training_ratio,
        bp_backprop_change[14],
        bp_weights_new[14]);

    backPropper_1 bp15(bp_dendrites[15],
        bp_weights[15],
        bp_axon,
        bp_backprop,
        bp_training_ratio,
        bp_backprop_change[15],
        bp_weights_new[15]);

    backPropper_1 bp16(bp_dendrites[16],
        bp_weights[16],
        bp_axon,
        bp_backprop,
        bp_training_ratio,
        bp_backprop_change[16],
        bp_weights_new[16]);

    backPropper_1 bp17(bp_dendrites[17],
        bp_weights[17],
        bp_axon,
        bp_backprop,
        bp_training_ratio,
        bp_backprop_change[17],
        bp_weights_new[17]);

    backPropper_1 bp18(bp_dendrites[18],
        bp_weights[18],
        bp_axon,
        bp_backprop,
        bp_training_ratio,
        bp_backprop_change[18],
        bp_weights_new[18]);

    backPropper_1 bp19(bp_dendrites[19],
        bp_weights[19],
        bp_axon,
        bp_backprop,
        bp_training_ratio,
        bp_backprop_change[19],
        bp_weights_new[19]);

    backPropper_1 bp20(bp_dendrites[20],
        bp_weights[20],
        bp_axon,
        bp_backprop,
        bp_training_ratio,
        bp_backprop_change[20],
        bp_weights_new[20]);

    backPropper_1 bp21(bp_dendrites[21],
        bp_weights[21],
        bp_axon,
        bp_backprop,
        bp_training_ratio,
        bp_backprop_change[21],
        bp_weights_new[21]);

    backPropper_1 bp22(bp_dendrites[22],
        bp_weights[22],
        bp_axon,
        bp_backprop,
        bp_training_ratio,
        bp_backprop_change[22],
        bp_weights_new[22]);

    backPropper_1 bp23(bp_dendrites[23],
        bp_weights[23],
        bp_axon,
        bp_backprop,
        bp_training_ratio,
        bp_backprop_change[23],
        bp_weights_new[23]);

    backPropper_1 bp24(bp_dendrites[24],
        bp_weights[24],
        bp_axon,
        bp_backprop,
        bp_training_ratio,
        bp_backprop_change[24],
        bp_weights_new[24]);

    backPropper_1 bp25(bp_dendrites[25],
        bp_weights[25],
        bp_axon,
        bp_backprop,
        bp_training_ratio,
        bp_backprop_change[25],
        bp_weights_new[25]);

    backPropper_1 bp26(bp_dendrites[26],
        bp_weights[26],
        bp_axon,
        bp_backprop,
        bp_training_ratio,
        bp_backprop_change[26],
        bp_weights_new[26]);

    backPropper_1 bp27(bp_dendrites[27],
        bp_weights[27],
        bp_axon,
        bp_backprop,
        bp_training_ratio,
        bp_backprop_change[27],
        bp_weights_new[27]);

    backPropper_1 bp28(bp_dendrites[28],
        bp_weights[28],
        bp_axon,
        bp_backprop,
        bp_training_ratio,
        bp_backprop_change[28],
        bp_weights_new[28]);

    backPropper_1 bp29(bp_dendrites[29],
        bp_weights[29],
        bp_axon,
        bp_backprop,
        bp_training_ratio,
        bp_backprop_change[29],
        bp_weights_new[29]);

    backPropper_1 bp30(bp_dendrites[30],
        bp_weights[30],
        bp_axon,
        bp_backprop,
        bp_training_ratio,
        bp_backprop_change[30],
        bp_weights_new[30]);

    backPropper_1 bp31(bp_dendrites[31],
        bp_weights[31],
        bp_axon,
        bp_backprop,
        bp_training_ratio,
        bp_backprop_change[31],
        bp_weights_new[31]);

    backPropper_t bpthresh(bp_weights[32],
        bp_backprop,
        bp_axon,
        bp_training_ratio,
        bp_weights_new[32]);

endmodule: backPropper

